library verilog;
use verilog.vl_types.all;
entity input_handler_tb is
end input_handler_tb;
