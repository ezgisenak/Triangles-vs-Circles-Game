/*module TrianglesVsCircles (
  input wire clk, 
  input wire reset,
  input wire logic_0_button,
  input wire logic_1_button,
  input wire activity_button,
  output wire vga_hsync,
  output wire vga_vsync,
  output wire [9:0] vga_red,
  output wire [9:0] vga_green,
  output wire [9:0] vga_blue
);

  // Game parameters
  parameter BOARD_SIZE = 10;
  parameter MAX_MOVES = 25;
  parameter WINNING_PLACEMENT = 4;
  
  typedef enum logic [2:0] {IDLE, TRIANGLES_TURN, CIRCLES_TURN, CHECK_WIN, GAME_OVER} state_t;
	state_t state, next_state;
	
	 typedef enum logic [1:0] {EMPTY = 2'b00, TRIANGLE = 2'b01, CIRCLE = 2'b10, OCCUPIED = 2'b11} piece_t;
	
  // Game state variables
  reg [1:0] board [0:BOARD_SIZE-1][0:BOARD_SIZE-1];
  reg current_player; // 0 for circle 1 for triangle
  reg [9:0] total_moves_triangles;
  reg [9:0] total_moves_circles;
  reg [9:0] recent_position_triangles;
  reg [9:0] recent_position_circles;
  reg [9:0] winning_placement_start_x;
  reg [9:0] winning_placement_start_y;
  reg [0:1] game_outcome;
  reg [3:0] move_counter;
  reg [9:0] erase_square_x;
  reg [9:0] erase_square_y;

  // VGA timing variables
  reg [10:0] hcount;
  reg [10:0] vcount;

  // Other internal signals
  wire [3:0] player_shape;
  
  // Game state initialization
  initial begin
    reset_game_state();
  end

  always_comb begin
    case(state)
      IDLE: begin
        // Idle state
      end
      TRIANGLES_TURN: begin
        // Triangles team's turn
      end
      CIRCLES_TURN: begin
        // Circles team's turn
      end
      CHECK_WIN: begin
        // Checking for a win
      end
      GAME_OVER: begin
        // Game over
      end
    endcase
  end
  
    always_ff @(posedge clk) begin
    if (reset) begin
      // reset logic
    end else if (logic_0_button) begin
      // add a '0' to the input buffer
    end else if (logic_1_button) begin
      // add a '1' to the input buffer
    end else if (activity_button) begin
      // interpret the input buffer as a move and make the move
    end
  end
	 
	   always_ff @(posedge clk) begin
    if (reset) begin
      // reset the display
    end else begin
      // update the display based on the game state
    end
  end
endmodule

  // Reset game state
  task reset_game_state;
    integer i, j;

    for (i = 0; i < BOARD_SIZE; i = i + 1) begin
      for (j = 0; j < BOARD_SIZE; j = j + 1) begin
        board[i][j] = 2'b00;
      end
	end
    endtask

	// Check if the move is valid
function automatic is_valid_move;
	
  input logic [3:0] x_input, // 4 bits for x coordinate
    input logic [3:0] y_input, // 4 bits for y coordinate

  // Check if the coordinates are within the board boundaries
 function logic is_valid_move(input [3:0] x, input [3:0] y);
    if(x >= SIZE || y >= SIZE || board[x][y] != EMPTY)
      return 0; // Invalid move
    else
      return 1; // Valid move
  endfunction
endfunction

endmodule
*/