/*module Display();

  // VGA timing generation
  always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
      hcount <= 0;
      vcount <= 0;
		state <= IDLE;
    end else if (vcount == 521 && hcount == 1280) begin
      state <= next_state;
		hcount <= 0;
      vcount <= 0;
    end else if (hcount == 1280) begin
		state <= next_state;
      hcount <= 0;
      vcount <= vcount + 1;
    end else begin
		state <= next_state;
      hcount <= hcount + 1;
    end
  end
  
  // VGA sync signals generation
  assign vga_hsync = (hcount >= 96 && hcount < 112) ? 1'b0 : 1'b1;
  assign vga_vsync = (vcount >= 2 && vcount < 34) ? 1'b0 : 1'b1;

  // VGA screen display generation
  always @(vcount, hcount) begin
    // VGA screen pixel generation logic
    // ...
    // Generate vga_red, vga_green, and vga_blue signals based on the current pixel

    // Update game state based on player inputs
		reg [3:0] x;
		
		always @* begin
		  if (activity_button) begin
			 x = {logic_1_button, logic_0_button};
		  end
		end
		  
      // Perform the move
      if (is_valid_move(x)) begin
        place_shape(x);
        update_game_state(x);
      end
    end
*/