library verilog;
use verilog.vl_types.all;
entity debounced_input_handler_tb is
end debounced_input_handler_tb;
